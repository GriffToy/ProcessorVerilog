// TCES 330, Spring 2016
// 5/28/2016
// Griffin Toyoda
// 16 bit 8-to-1 mux

module Mux16w_8to1(S, Q, R, T, U, V, W, X, Y, M);
	input [15:0] Q, R, T, U, V, W, X, Y;	// Input lines
	input [2:0] S;				            // Selection lines
	output [15:0] M;

	wire A, B, C;

	Mux8_1 u1(Q[0], R[0], T[0], U[0], V[0], W[0], X[0], Y[0], S, M[0]);
	Mux8_1 u2(Q[1], R[1], T[1], U[1], V[1], W[1], X[1], Y[1], S, M[1]);
	Mux8_1 u3(Q[2], R[2], T[2], U[2], V[2], W[2], X[2], Y[2], S, M[2]);
	Mux8_1 u4(Q[3], R[3], T[3], U[3], V[3], W[3], X[3], Y[3], S, M[3]);
	Mux8_1 u5(Q[4], R[4], T[4], U[4], V[4], W[4], X[4], Y[4], S, M[4]);
	Mux8_1 u6(Q[5], R[5], T[5], U[5], V[5], W[5], X[5], Y[5], S, M[5]);
	Mux8_1 u7(Q[6], R[6], T[6], U[6], V[6], W[6], X[6], Y[6], S, M[6]);
	Mux8_1 u8(Q[7], R[7], T[7], U[7], V[7], W[7], X[7], Y[7], S, M[7]);
	Mux8_1 u9(Q[8], R[8], T[8], U[8], V[8], W[8], X[8], Y[8], S, M[8]);
	Mux8_1 u10(Q[9], R[9], T[9], U[9], V[9], W[9], X[9], Y[9], S, M[9]);
	Mux8_1 u11(Q[10], R[10], T[10], U[10], V[10], W[10], X[10], Y[10], S, M[10]);
	Mux8_1 u12(Q[11], R[11], T[11], U[11], V[11], W[11], X[11], Y[11], S, M[11]);
	Mux8_1 u13(Q[12], R[12], T[12], U[12], V[12], W[12], X[12], Y[12], S, M[12]);
	Mux8_1 u14(Q[13], R[13], T[13], U[13], V[13], W[13], X[13], Y[13], S, M[13]);
	Mux8_1 u15(Q[14], R[14], T[14], U[14], V[14], W[14], X[14], Y[14], S, M[14]);
	Mux8_1 u16(Q[15], R[15], T[15], U[15], V[15], W[15], X[15], Y[15], S, M[15]);
	
endmodule